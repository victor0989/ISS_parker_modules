module ROM_MEMORY (
    input  [35:0] addr,
    output reg [63:0] data_val
);

    always @* begin
        case (addr[35:3]) // Ignorar los 3 bits menos significativos
            33'h20000000: data_val = 64'h1400004f_040000ff;
            33'h20000001: data_val = 64'h17000a01_1900474e;
            33'h20000002: data_val = 64'h17003a41_00380180;
            33'h20000003: data_val = 64'h1900638e_03000037;
            33'h20000004: data_val = 64'h1900630e_00010731;
            33'h20000005: data_val = 64'h14ffffc8_04ff6088;
            33'h20000006: data_val = 64'h13001810_17003381;
            33'h20000007: data_val = 64'h1900448e_19fffc40;
            33'h20000008: data_val = 64'h03000074_03000035;
            33'h20000009: data_val = 64'h03000037_04000006;
            33'h2000000A: data_val = 64'h19005d8e_1f000150;
            33'h2000000B: data_val = 64'h01000155_01ffff44;
            33'h2000000C: data_val = 64'h12fff400_19005c4e;
            33'h2000000D: data_val = 64'h25000160_10001060;
            33'h2000000E: data_val = 64'h17002d11_190040ce;
            33'h2000000F: data_val = 64'h19fff880_17002aa1;
            33'h20000010: data_val = 64'h1900400e_15636f01;
            33'h20000011: data_val = 64'h166c6411_16626f11;
            33'h20000012: data_val = 64'h046f7411_14000042;
            33'h20000013: data_val = 64'h04000022_04000003;
            33'h20000014: data_val = 64'h04000004_1a000070;
            33'h20000015: data_val = 64'h0a2a2a2a_2a2a2042;
            33'h20000016: data_val = 64'h4f4f5420_50524f47;
            33'h20000017: data_val = 64'h52414d20_284d4242;
            33'h20000018: data_val = 64'h6f6f7465_722e7329;
            33'h20000019: data_val = 64'h202a2a2a_2a2a0a20;
            33'h2000001A: data_val = 64'h2020456e_74657220;
            33'h2000001B: data_val = 64'h64617461_20696e20;
            33'h2000001C: data_val = 64'h74686973_20666f72;
            33'h2000001D: data_val = 64'h6d61743a_0a202020;
            33'h2000001E: data_val = 64'h20203820_62797465;
            33'h2000001F: data_val = 64'h733a204e_3d6e756d;
            33'h20000020: data_val = 64'h62657220_6f662064;
            33'h20000021: data_val = 64'h61746120_62797465;
            33'h20000022: data_val = 64'h730a2020_20202038;
            33'h20000023: data_val = 64'h20627974_65733a20;
            33'h20000024: data_val = 64'h413d6164_64726573;
            33'h20000025: data_val = 64'h73206174_20776869;
            33'h20000026: data_val = 64'h63682074_6f20706c;
            33'h20000027: data_val = 64'h61636520_74686520;
            33'h20000028: data_val = 64'h64617461_20627974;
            33'h20000029: data_val = 64'h65732028_6e6f726d;
            33'h2000002A: data_val = 64'h616c6c79_20303030;
            33'h2000002B: data_val = 64'h30303030_30303030;
            33'h2000002C: data_val = 64'h30303030_38290a20;
            33'h2000002D: data_val = 64'h20202020_4e206279;
            default: data_val = 64'h00000000_00000000;
        endcase
    end
endmodule // ROM_MEMORY

